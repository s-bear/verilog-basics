`timescale 1ns/10ps

/*
test_debounce.v
2019-04-11 Samuel B Powell
samuel.powell@uq.edu.au

*/


module test_debounce;
initial begin
    $dumpfile("test_debounce.fst");
    $dumpvars(-1,test_debounce);
end



endmodule